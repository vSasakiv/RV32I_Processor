module template (
  ports
);
  
endmodule