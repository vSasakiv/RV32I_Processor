module test #(
  parameters
) (
  initial begin
    $display("Test")
  end
);

endmodule