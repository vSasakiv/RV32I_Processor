module template #(
  parameters
) (
  ports
);

endmodule