module cpu #(

) (

);

endmodule