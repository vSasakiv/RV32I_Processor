module cpu_mod #(
  parameters
) (
  ports
);
  
endmodule